// =============================================================================
// MAZE网络QoS仲裁器模块
// =============================================================================
// 功能说明：
// 1. 基于QoS优先级的固定优先级仲裁器
// 2. 默认支持4个请求输入的仲裁，可通过配置WIDTH实现任意输入
// 3. 高QoS请求具有绝对优先权
// 4. 相同QoS级别时采用固定优先级仲裁
// 5. 组合逻辑实现，1个时钟周期完成仲裁
// =============================================================================

module arbiter #(
    parameter WIDTH = 4                    // 仲裁器输入宽度，默认4个输入
) (
    // 仲裁器输入接口
    input  logic [WIDTH-1:0] req,          // 请求信号，1表示有请求
    input  logic [WIDTH-1:0] qos,          // QoS优先级信号，1表示高优先级

    // 仲裁器输出接口
    output logic [WIDTH-1:0] gnt           // 授权信号，1表示获得授权
);

// =============================================================================
// QoS仲裁逻辑实现
// =============================================================================
// 仲裁策略：
// 1. 如果有高QoS请求(qos=1)，则优先处理高QoS请求
// 2. 高QoS请求中采用最低位的固定优先级
// 3. 如果没有高QoS请求，则处理普通请求(req=1)
// 4. 普通请求中采用最低位的固定优先级
// 5. 使用位操作实现高效的优先级编码
// =============================================================================

assign gnt = (|qos) ? (qos & (~(qos-1))) : (req & (~(req-1)));

endmodule
