interface pkt_con_if;
   

endinterface : pkt_con_if